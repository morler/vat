module printer

const buf_size = 64 * 1024

pub interface Printer {
	print()
}
